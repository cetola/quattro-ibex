package vip_pkg;

`include "coverage.svh"
`include "tester.svh"
`include "scoreboard.svh"
`include "testbench.svh"

endpackage : vip_pkg
